
module top (
    output  logic[7:0]      led
);

    assign led = 8'hf3;

    system system_i ();
    
endmodule

